module controller (
    input logic clk,
    output logic load_sreg,
    output logic transmit_pixel,
    output logic
);

endmodule
